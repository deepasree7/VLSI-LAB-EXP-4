module T_flipflop(t,clk,rstn,q);
input t,clk,rstn;
output reg q;
always @(posedge clk) begin
if (!rstn)
q<=0;
else
if (t)
q<= ~q;
else
q<= q;
end
endmodule
